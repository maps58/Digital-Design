{\rtf1\ansi\ansicpg1252\deff0\deflang2058{\fonttbl{\f0\fnil\fcharset0 Calibri;}}
{\*\generator Msftedit 5.41.21.2510;}\viewkind4\uc1\pard\sl240\slmult1\lang10\f0\fs28\par
library IEEE;\par
use IEEE.STD_LOGIC_1164.ALL;\par
\par
entity decode_2to4_top is\par
    Port ( sw : in  STD_LOGIC_VECTOR (2 downto 0);  -- 2-bit input\par
               led : out STD_LOGIC_VECTOR (3 downto 0);  -- 4-bit output\par
              \par
end decode_2to4_top;\par
\par
architecture Behavioral of decode_2to4_top is\par
signal a: std_ logic _vector (1 downto 0);\par
signal en: std_logic;\par
signal x: std_logic_vector (3 downto 0);\par
begin\par
process (A, EN)\par
begin\par
    X <= "1111";        -- default output value\par
    if (EN = '1') then  -- active high enable pin\par
        case A is\par
            when "00" => X(0) <= '0';\par
            when "01" => X(1) <= '0';\par
            when "10" => X(2) <= '0';\par
            when "11" => X(3) <= '0';\par
            when others => X <= "1111";\par
        end case;\par
    end if;\par
end process;\par
\par
led <= x(3 downto 0);\par
a<= sw(1 downto 0);\par
en<= sw(2);\par
\par
\par
end Behavioral;\par
}
 