{\rtf1\ansi\ansicpg1252\deff0\deflang2058{\fonttbl{\f0\fnil\fcharset0 Calibri;}{\f1\fnil\fcharset0 Courier New;}}
{\*\generator Msftedit 5.41.21.2510;}\viewkind4\uc1\pard\sl276\slmult1\qc\lang10\f0\fs36 PRACTICA 9: CONTADORES SINCRONOS Y ASINCRONOS (Contador de decada_comportamental)\par
\pard\sl276\slmult1\par
\par
\pard\lang2058\f1\fs28 library ieee;\par
use ieee.std_logic_1164.all;\par
use ieee.std_logic_unsigned.all;\par
\tab  \par
entity contador is port(\par
clk, reset:in std_logic;\par
conta: out std_logic_vector(3 downto 0));\par
end contador; \tab  \par
\tab  \par
\tab  \par
architecture archicontador of contador is\par
signal temp: std_logic_vector (3 downto 0);\par
begin\par
process (clk,reset)\par
begin\par
  if reset = '1' then\par
     temp <= "0000";\par
        elsif (clk'event and clk= '1') then\par
\tab\tab   \par
\tab\tab   \par
\tab\tab      if  temp = "1001" then\par
\tab\tab\tab    temp <="0000" ;\par
\tab\tab\tab\tab else\par
         \tab\tab\par
\tab\tab\tab temp <= temp + 1;\par
         \tab\tab\par
\tab\tab   \par
\tab   end if;\par
  end if;\par
end process;\par
conta <= temp;\par
end archicontador;\par
\pard\sl276\slmult1\lang10\f0\fs36\par
}
 