library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Numeric_Std.all;

entity GrayCounter3p_tb is
end;

architecture bench of GrayCounter3p_tb is

  component GrayCounter3p
          Port ( rst : in  STD_LOGIC;
          clk : in  STD_LOGIC;
  	      sel : in  STD_LOGIC;
          GrayCount : out  STD_LOGIC_VECTOR(2 downto 0));
  end component;

  signal rst: STD_LOGIC;
  signal clk: STD_LOGIC;
  signal sel: STD_LOGIC;
  signal GrayCount: STD_LOGIC_VECTOR(2 downto 0);

  constant clock_period: time := 10 ns;
  signal stop_the_clock: boolean;

begin

  uut: GrayCounter3p port map ( rst=> rst,clk=> clk,sel=> sel,GrayCount => GrayCount );

  stimulus: process
  begin

  rst <= '0'; sel <='0'; wait for 50 ns;
  rst <= '1'; sel <= '1'; wait for 700 ns;
  sel <= '0'; wait for 200 ns;
  rst <= '0'; wait for 100 ns;

 end process;
 
 clocking: process
  begin
    while not stop_the_clock loop
      clk <= '0', '1' after clock_period / 2;
      wait for clock_period;
    end loop;
    wait;
  end process;
end;
