{\rtf1\ansi\ansicpg1252\deff0\deflang2058{\fonttbl{\f0\fnil\fcharset0 Calibri;}}
{\*\generator Msftedit 5.41.21.2510;}\viewkind4\uc1\pard\sl276\slmult1\qc\lang10\b\f0\fs28 PRACTICA 10: REGISTROS (PIPO_ COMPORTAMENTAL)\par
\pard\sl276\slmult1\b0\fs22\par
\fs32 library ieee;  \par
use ieee.std_logic_1164.all;  \par
 \par
entity flop is  \par
  port(CLK, CE, PRE : in std_logic;  \par
        D : in  std_logic_vector (3 downto 0);  \par
        Q : out std_logic_vector (3 downto 0));  \par
end flop; \par
architecture archi of flop is  \par
  begin  \par
    process (CLK, PRE)  \par
      begin  \par
        if (PRE='1') then  \par
          Q <= "1111";  \par
        elsif (CLK'event and CLK='1')then  \par
          if (CE='1') then  \par
            Q <= D;  \par
          end if;  \par
        end if;  \par
    end process;  \par
end archi; \par
}
 